----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:    13:36:12 12/09/2018
-- Design Name:
-- Module Name:    gray_counter - Behavioral
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

--! @brief Entity for a 4-bit Gray code counter.
--!
--! This entity implements a 4-bit Gray code counter with output to a 7-segment
--! display. The counter is controlled by a push button and a clock signal.
entity gray_counter is
    Port (
        --! @brief Push button input to enable/disable counting.
        --!
        --! When '1', the counter advances through the Gray code sequence.
        --! When '0', the counter is paused.
        pb : in STD_LOGIC;
        --! @brief System clock input.
        clk : in  STD_LOGIC;
        --! @brief 4-bit output to control the 7-segment display anodes.
        en : out  STD_LOGIC_VECTOR (3 downto 0);
        --! @brief 8-bit output for the 7-segment display segments.
        led : out  STD_LOGIC_VECTOR (7 downto 0)
    );
end gray_counter;

architecture Behavioral of gray_counter is
    --! @brief Stores the current 4-bit Gray code value.
    signal tmp: STD_LOGIC_VECTOR (3 downto 0):= "0000";
    --! @brief Slow clock signal generated by a clock divider.
    signal my_clk: STD_LOGIC;
    --! @brief 4-bit signal to select which 7-segment display is active.
    signal sel: unsigned (3 downto 0) := "1110";
    --! @brief 8-bit signal to control the segments of the 7-segment display.
    signal tmpLED: unsigned (7 downto 0) := "00000000";
begin

    -- Assign internal signals to output ports
    en <= std_logic_vector(sel);
    led <= std_logic_vector(tmpLED);

    --! @brief Process to drive the 7-segment display.
    --!
    --! This process determines which segments to light up based on the
    --! current Gray code value (tmp) and the active display (sel).
    --! When pb is '1', it displays '0' or '1'.
    --! When pb is '0', it displays characters 's', 'a', 'p'.
    process(sel, pb, tmp)
    begin
        if(pb = '1') then
            case sel is
            when "1110" =>
                if tmp(0) = '0' then
                    tmpLED <= x"c0"; -- '0'
                else
                    tmpLED <= x"f9"; -- '1'
                end if;
            when "1101" =>
                if tmp(1) = '0' then
                    tmpLED <= x"c0"; -- '0'
                else
                    tmpLED <= x"f9"; -- '1'
                end if;
            when "1011" =>
                if tmp(2) = '0' then
                    tmpLED <= x"c0"; -- '0'
                else
                    tmpLED<= x"f9"; -- '1'
                end if;
            when "0111" =>
                if tmp(3) = '0' then
                    tmpLED <= x"c0"; -- '0'
                else
                    tmpLED <= x"f9"; -- '1'
                end if;
            when others =>
                tmpLED <= (others => '0');
            end case;
        else
            case sel is
            when "1110" =>
                if tmp(0) = '0' then
                    tmpLED <= x"92"; -- 's'
                end if;
            when "1101" =>
                if tmp(1) = '0' then
                    tmpLED <= x"92"; -- 's'
                end if;
            when "1011" =>
                if tmp(2) = '0' then
                    tmpLED <= x"88"; -- 'a'
                end if;
            when "0111" =>
                if tmp(3) = '0' then
                    tmpLED <= x"8c"; -- 'p'
                end if;
            when others =>
                tmpLED <= (others => '0');
            end case;
        end if;
    end process;

    --! @brief Process to rotate the 7-segment display selection.
    --!
    --! This process creates a scanning effect for the 4-digit 7-segment
    --! display by rotating the 'sel' signal.
    process(clk)
        variable counter : integer range 0 to 5000 := 0;
    begin
        if(rising_edge(clk)) then
            counter := counter + 1;
            if counter = 2499 then
                counter := 0;
                sel <= sel ror 1;
            end if;
        end if;
    end process;

    --! @brief Process to generate a slow clock signal (my_clk).
    --!
    --! This process divides the main clock 'clk' to create a slower clock
    --! 'my_clk' that controls the Gray code counter's update rate.
    process(clk)
        variable cc : integer range 0 to 12000000 := 0;
    begin
        if(rising_edge(clk)) then
            cc := cc + 1;
            if(cc = 11999999) then
                cc := 0;
                my_clk <= not my_clk;
            end if;
        end if;
    end process;

    --! @brief Process to generate the 4-bit Gray code sequence.
    --!
    --! This process updates the Gray code value 'tmp' on the rising edge of
    --! 'my_clk' only when the push button 'pb' is pressed.
    process(my_clk)
    begin
        if(rising_edge(my_clk)) then
            if(pb = '1') then
                case tmp is
                    when "0000" => tmp <= "0001";
                    when "0001" => tmp <= "0011";
                    when "0011" => tmp <= "0010";
                    when "0010" => tmp <= "0110";
                    when "0110" => tmp <= "0111";
                    when "0111" => tmp <= "0101";
                    when "0101" => tmp <= "0100";
                    when "0100" => tmp <= "1100";
                    when "1100" => tmp <= "1101";
                    when "1101" => tmp <= "1111";
                    when "1111" => tmp <= "1110";
                    when "1110" => tmp <= "1010";
                    when "1010" => tmp <= "1011";
                    when "1011" => tmp <= "1001";
                    when "1001" => tmp <= "1000";
                    when "1000" => tmp <= "0000";
                    when others => tmp <= "0000";
                end case;
            end if;
        end if;
    end process;

end Behavioral;
